(** Coq module loading the different ML components of the plugin **)

Declare ML Module "error".
Declare ML Module "modules".
Declare ML Module "libraries".
Declare ML Module "commands".

