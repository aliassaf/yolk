(** Coq module loading the Yolk plugin **)

Declare ML Module "yolk_plugin".

