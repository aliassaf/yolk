(** Coq module loading the different ML components of the plugin **)

Declare ML Module "error".
Declare ML Module "export".
Declare ML Module "commands".

